layer;name=initialization;
entity;name=MainController;layer=initialization
component;name=CreateSpheres;prefix=gameplay/spherebuilder;entity=MainController