layer;name=initialization;
entity;name=MainController;layer=initialization
component;name=TargetPractice;prefix=gameplay/targetPractice;entity=MainController